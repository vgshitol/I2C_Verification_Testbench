package wb_pkg;

  import ncsu_pkg::*;

  `include "ncsu_macros.svh"
  `include "src/wb_header.svh"
  `include "src/wb_configuration.svh"
  `include "src/wb_transaction.svh"
  `include "src/wb_transaction_random.svh"
  `include "src/wb_driver.svh"
  `include "src/wb_monitor.svh"
  `include "src/wb_coverage.svh"
  `include "src/wb_agent.svh"

endpackage




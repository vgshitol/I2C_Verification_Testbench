package wb_pkg;

  `include "src/wb_configuration.svh"
  `include "src/wb_agent.svh"
  `include "src/wb_driver.svh"
  `include "src/wb_monitor.svh"
  `include "src/wb_transaction.svh"
 
endpackage
